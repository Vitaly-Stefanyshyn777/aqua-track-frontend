<svg xmlns="http://www.w3.org/2000/svg" aria-hidden="true" style="position:absolute;width:0;height:0;overflow:hidden">
  <defs>
    <symbol id="icon-edit-2" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3.6" d="M22.666 4a3.766 3.766 0 0 1 4.109-.817 3.781 3.781 0 0 1 2.041 2.04 3.764 3.764 0 0 1 0 2.886 3.756 3.756 0 0 1-.817 1.223l-18 18-7.333 2 2-7.333 18-18z"/>
    </symbol>
    <symbol id="icon-emojione-v1_white-exclamation-mark" viewBox="0 0 32 32">
      <path fill="#9be1a0" d="M13.474 18.545c.121 1.266.328 2.206.611 2.827.287.618.796.927 1.532.927.137 0 .261-.022.383-.047.125.025.247.047.386.047.734 0 1.244-.308 1.53-.927.285-.62.488-1.561.611-2.827l.653-9.771c.122-1.905.184-3.271.184-4.101 0-1.129-.295-2.01-.886-2.643-.593-.632-1.372-.948-2.337-.948-.052 0-.09.012-.14.014-.048-.002-.087-.014-.137-.014-.967 0-1.745.316-2.337.948s-.888 1.515-.888 2.643c0 .83.06 2.196.184 4.101l.652 9.77zm2.551 7.325c-.937 0-1.733.295-2.394.886s-.992 1.31-.992 2.153c0 .951.335 1.701 1 2.244.668.544 1.447.816 2.338.816.906 0 1.697-.268 2.373-.806.675-.536 1.012-1.289 1.012-2.254 0-.843-.323-1.561-.969-2.153s-1.436-.887-2.37-.887z" style="fill:var(--color1, #9be1a0)"/>
    </symbol>
    <symbol id="icon-Ellipse-2" viewBox="0 0 35 32">
      <path fill="#fff" stroke="#9be1a0" stroke-width="2.667" d="M32 16c0 8.1-6.566 14.667-14.667 14.667S2.666 24.101 2.666 16c0-8.1 6.566-14.667 14.667-14.667S32 7.899 32 16z" style="fill:var(--color1, #fff);stroke:var(--color2, #9be1a0)"/>
    </symbol>
    <symbol id="icon-eye" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="2.88" d="M1.333 16S6.666 5.333 16 5.333 30.667 16 30.667 16 25.334 26.667 16 26.667 1.333 16 1.333 16z"/>
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="2.88" d="M16 20a4 4 0 1 0 0-8 4 4 0 0 0 0 8z"/>
    </symbol>
    <symbol id="icon-eye-off" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="2.88" d="M23.92 23.92A13.43 13.43 0 0 1 16 26.667C6.667 26.667 1.333 16 1.333 16A24.605 24.605 0 0 1 8.08 8.08m5.12-2.427a12.161 12.161 0 0 1 2.8-.32C25.333 5.333 30.667 16 30.667 16a24.646 24.646 0 0 1-2.88 4.253m-8.961-1.426a4.01 4.01 0 0 1-2.855 1.273 3.978 3.978 0 0 1-1.569-.291 3.984 3.984 0 0 1-2.21-2.21 3.995 3.995 0 0 1 .983-4.424M1.333 1.333l29.333 29.333"/>
    </symbol>
    <symbol id="icon-log-out" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3" d="M12 28H6.667A2.668 2.668 0 0 1 4 25.333V6.666a2.668 2.668 0 0 1 2.667-2.667H12M21.334 22.667 28.001 16l-6.667-6.667M28 16H12"/>
    </symbol>
    <symbol id="icon-mage_water-glass-fill" viewBox="0 0 31 32">
      <path fill="#9be1a0" d="M26.955 5.226c-.095-.321-.254-.616-.468-.868s-.477-.452-.772-.589a2.087 2.087 0 0 0-.937-.21H6.562a1.83 1.83 0 0 0-.937.197c-.301.139-.57.345-.785.604a2.36 2.36 0 0 0-.468.866 2.392 2.392 0 0 0-.089.984l2.076 18.377a5.202 5.202 0 0 0 1.633 3.255 4.78 4.78 0 0 0 3.253 1.313h8.861a4.804 4.804 0 0 0 3.266-1.313 5.316 5.316 0 0 0 1.62-3.255l1.127-10.331v-.158l.873-7.876a2.724 2.724 0 0 0-.038-.998zM14.17 25.375h-1.266a3.573 3.573 0 0 1-2.215-.945 3.744 3.744 0 0 1-1.139-2.192l-.304-2.258c-.039-.344.053-.691.258-.965s.504-.455.835-.503.667.04.936.246.45.512.503.854l.304 2.232c.034.244.151.467.329.63a1 1 0 0 0 .646.276h1.266c.336 0 .658.138.895.384s.371.58.371.928-.133.682-.371.928a1.242 1.242 0 0 1-.895.384h-.152zm10.127-12.116c-2.671.538-4.949.643-7.367-1.313-3-2.455-6.633-1.667-10.127-.381L6.17 5.999a.41.41 0 0 1 0-.171.337.337 0 0 1 .089-.144.257.257 0 0 1 .127-.105.262.262 0 0 1 .152 0h18.38a.53.53 0 0 1 .127.105.314.314 0 0 1 .076.144.304.304 0 0 1 0 .184l-.823 7.246z" style="fill:var(--color1, #9be1a0)"/>
    </symbol>
    <symbol id="icon-pie-chart-02" viewBox="0 0 32 32">
      <path fill="none" stroke="#323f47" stroke-linecap="round" stroke-linejoin="round" stroke-width="2.667" d="M22.933 18.667c.369 0 .554 0 .704.082a.713.713 0 0 1 .293.324c.067.157.05.324.016.659a10.665 10.665 0 0 1-12.694 9.397c-2.069-.412-3.97-1.428-5.462-2.919s-2.508-3.392-2.919-5.461a10.666 10.666 0 0 1 9.397-12.694c.334-.034.502-.05.659.016.13.055.257.17.324.293.082.15.082.334.082.704v8.533c0 .373 0 .56.073.703a.67.67 0 0 0 .291.291c.143.073.329.073.703.073h8.533z" style="stroke:var(--color2, #323f47)"/>
      <path fill="none" stroke="#9be1a0" stroke-linecap="round" stroke-linejoin="round" stroke-width="2.667" d="M18.667 3.733c0-.369 0-.554.082-.704a.713.713 0 0 1 .324-.293c.157-.067.324-.05.659-.016a10.67 10.67 0 0 1 9.549 9.549c.033.334.05.502-.016.659a.704.704 0 0 1-.293.324c-.15.082-.334.082-.704.082h-8.533c-.373 0-.56 0-.703-.073a.67.67 0 0 1-.291-.291c-.073-.143-.073-.329-.073-.703V3.734z" style="stroke:var(--color1, #9be1a0)"/>
    </symbol>
    <symbol id="icon-minus1" viewBox="0 0 32 32">
      <path stroke-width="1.116" d="M16 .558C24.528.558 31.442 7.472 31.442 16S24.528 31.442 16 31.442.558 24.528.558 16 7.472.558 16 .558z"/>
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="1.339" d="M10.286 16h11.429"/>
    </symbol>
    <symbol id="icon-plus" viewBox="0 0 32 32">
      <path stroke-linejoin="round" stroke-linecap="round" stroke-miterlimit="4" stroke-width="3" d="M16 6.667v18.667"></path>
      <path stroke-linejoin="round" stroke-linecap="round" stroke-miterlimit="4" stroke-width="3" d="M6.667 16h18.667"></path>
    </symbol>
    <symbol id="icon-plus2" viewBox="0 0 32 32">
      <path stroke-width="1.116" d="M16 .558C24.528.558 31.442 7.472 31.442 16S24.528 31.442 16 31.442.558 24.528.558 16 7.472.558 16 .558z"/>
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="1.339" d="M16 10.286v11.429M10.286 16h11.429"/>
    </symbol>
    <symbol id="icon-settings" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3" d="M16 20a4 4 0 1 0 0-8 4 4 0 0 0 0 8z"/>
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3" d="M25.867 20a2.205 2.205 0 0 0 .44 2.427l.08.08a2.672 2.672 0 0 1 .782 1.886 2.672 2.672 0 0 1-1.648 2.465 2.672 2.672 0 0 1-2.907-.579l-.08-.08a2.197 2.197 0 0 0-2.427-.44 2.2 2.2 0 0 0-1.334 2.013v.227a2.668 2.668 0 0 1-5.334 0v-.12a2.196 2.196 0 0 0-1.44-2.013 2.205 2.205 0 0 0-2.427.44l-.08.08a2.672 2.672 0 0 1-1.886.782 2.672 2.672 0 0 1-2.465-1.648 2.672 2.672 0 0 1 .579-2.907l.08-.08a2.197 2.197 0 0 0 .44-2.427 2.2 2.2 0 0 0-2.013-1.334H4a2.668 2.668 0 0 1 0-5.334h.12a2.196 2.196 0 0 0 2.013-1.44 2.2 2.2 0 0 0-.44-2.427l-.08-.08a2.666 2.666 0 0 1 .865-4.352 2.668 2.668 0 0 1 2.908.579l.08.08a2.197 2.197 0 0 0 2.427.44H12a2.2 2.2 0 0 0 1.334-2.013v-.227a2.668 2.668 0 0 1 5.334 0v.12a2.203 2.203 0 0 0 1.334 2.013 2.208 2.208 0 0 0 2.427-.44l.08-.08a2.672 2.672 0 0 1 1.886-.782 2.672 2.672 0 0 1 2.465 1.647 2.668 2.668 0 0 1-.579 2.907l-.08.08a2.197 2.197 0 0 0-.44 2.427v.107a2.2 2.2 0 0 0 2.013 1.334h.227a2.668 2.668 0 0 1 0 5.334h-.12a2.203 2.203 0 0 0-2.013 1.334z"/>
    </symbol>
    <symbol id="icon-down" viewBox="0 0 32 32">
      <path stroke-linejoin="round" stroke-linecap="round" stroke-miterlimit="4" stroke-width="3" d="M8 12l8 8 8-8"></path>
    </symbol>
    <symbol id="icon-trash-04" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3" d="M12 4h8"/>
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3.6" d="M4 8h24m-2.667 0-.935 14.026c-.14 2.104-.21 3.156-.665 3.954a4.007 4.007 0 0 1-1.731 1.62c-.826.4-1.881.4-3.99.4h-4.025c-2.109 0-3.163 0-3.99-.4a4.001 4.001 0 0 1-1.731-1.62c-.455-.798-.525-1.85-.665-3.954L6.666 8"/>
    </symbol>
    <symbol id="icon-upload" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="2.88" d="M28 20v5.333A2.668 2.668 0 0 1 25.333 28H6.666a2.668 2.668 0 0 1-2.667-2.667V20M22.666 10.667 15.999 4l-6.667 6.667M16 4v16"/>
    </symbol>
    <symbol id="icon-x-1" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3.429" d="M24 8 8 24M8 8l16 16"/>
    </symbol>
    <symbol id="icon-google-icon" viewBox="0 0 32 32">
<path fill="#fbbc05" style="fill: var(--color1, #fbbc05)" d="M6.885 16c0-1.016 0.169-1.99 0.47-2.904l-5.273-4.026c-1.028 2.086-1.607 4.437-1.607 6.93 0 2.491 0.578 4.841 1.604 6.925l5.27-4.034c-0.298-0.91-0.465-1.88-0.465-2.891z"></path>
<path fill="#eb4335" style="fill: var(--color2, #eb4335)" d="M16.142 6.756c2.208 0 4.201 0.782 5.768 2.062l4.558-4.551c-2.777-2.418-6.338-3.911-10.326-3.911-6.191 0-11.512 3.541-14.060 8.714l5.273 4.026c1.215-3.688 4.678-6.34 8.788-6.34z"></path>
<path fill="#34a853" style="fill: var(--color3, #34a853)" d="M16.142 25.244c-4.11 0-7.573-2.652-8.788-6.34l-5.273 4.026c2.548 5.174 7.869 8.715 14.060 8.715 3.821 0 7.469-1.357 10.208-3.899l-5.005-3.869c-1.412 0.89-3.19 1.368-5.203 1.368z"></path>
<path fill="#4285f4" style="fill: var(--color4, #4285f4)" d="M31.097 16c0-0.924-0.142-1.92-0.356-2.844h-14.598v6.044h8.403c-0.42 2.061-1.564 3.645-3.2 4.676l5.005 3.869c2.876-2.669 4.747-6.646 4.747-11.745z"></path>
</symbol>

  </defs>
</svg>

<!-- GPT написало які іконки використовуються нище для зручності, якщо не зрозуміло підключіть самостійно -->

<!-- 
<svg xmlns="http://www.w3.org/2000/svg" aria-hidden="true" style="position:absolute;width:0;height:0;overflow:hidden">
  <defs>

    <!-- Іконка редагування (олівець), зазвичай використовується для кнопки "Редагувати" -->
    <symbol id="icon-edit-2" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3.6"
            d="M22.666 4a3.766 3.766 0 0 1 4.109-.817 3.781 3.781 0 0 1 2.041 2.04 
               3.764 3.764 0 0 1 0 2.886 3.756 3.756 0 0 1-.817 1.223l-18 18-7.333 2 2-7.333 18-18z"/>
    </symbol>

    <!-- Білий знак оклику, використовується для попереджень або сповіщень -->
    <symbol id="icon-emojione-v1_white-exclamation-mark" viewBox="0 0 32 32">
      <path fill="#9be1a0"
            d="M13.474 18.545c.121 1.266.328 2.206.611 2.827.287.618.796.927 1.532.927.137 0 .261-.022.383-.047 
               .125.025.247.047.386.047.734 0 1.244-.308 1.53-.927.285-.62.488-1.561.611-2.827l.653-9.771c.122-1.905.184-3.271.184-4.101 
               0-1.129-.295-2.01-.886-2.643-.593-.632-1.372-.948-2.337-.948-.052 0-.09.012-.14.014-.048-.002-.087-.014-.137-.014-.967 0 
               -1.745.316-2.337.948s-.888 1.515-.888 2.643c0 .83.06 2.196.184 4.101l.652 9.77z"/>
    </symbol>

    <!-- Коло (еліпс), може бути використане як індикатор статусу -->
    <symbol id="icon-Ellipse-2" viewBox="0 0 35 32">
      <path fill="#fff" stroke="#9be1a0" stroke-width="2.667"
            d="M32 16c0 8.1-6.566 14.667-14.667 14.667S2.666 24.101 2.666 16c0-8.1 6.566-14.667 14.667-14.667S32 7.899 32 16z"/>
    </symbol>

    <!-- Іконка "Око" - використовується для показу пароля або попереднього перегляду контенту -->
    <symbol id="icon-eye" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="2.88"
            d="M1.333 16S6.666 5.333 16 5.333 30.667 16 30.667 16 25.334 26.667 16 26.667 1.333 16 1.333 16z"/>
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="2.88"
            d="M16 20a4 4 0 1 0 0-8 4 4 0 0 0 0 8z"/>
    </symbol>

    <!-- Іконка "Око закрите" (перекреслене око) - використовується для приховування пароля -->
    <symbol id="icon-eye-off" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="2.88"
            d="M23.92 23.92A13.43 13.43 0 0 1 16 26.667C6.667 26.667 1.333 16 1.333 16 
               A24.605 24.605 0 0 1 8.08 8.08m5.12-2.427a12.161 12.161 0 0 1 2.8-.32C25.333 5.333 30.667 16 
               30.667 16a24.646 24.646 0 0 1-2.88 4.253"/>
    </symbol>

    <!-- Іконка "Вихід" - використовується для кнопки "Вийти" -->
    <symbol id="icon-log-out" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3"
            d="M12 28H6.667A2.668 2.668 0 0 1 4 25.333V6.666a2.668 2.668 0 0 1 2.667-2.667H12M21.334 22.667 28.001 16l-6.667-6.667M28 16H12"/>
    </symbol>

    <!-- Іконка "Склянка з водою" - використовується для відстеження гідратації -->
    <symbol id="icon-mage_water-glass-fill" viewBox="0 0 31 32">
      <path fill="#9be1a0"
            d="M26.955 5.226c-.095-.321-.254-.616-.468-.868s-.477-.452-.772-.589a2.087 2.087 0 0 0-.937-.21H6.562a1.83 
               1.83 0 0 0-.937.197c-.301.139-.57.345-.785.604a2.36 2.36 0 0 0-.468.866 2.392 2.392 0 0 0-.089.984l2.076 
               18.377a5.202 5.202 0 0 0 1.633 3.255 4.78 4.78 0 0 0 3.253 1.313h8.861a4.804 4.804 0 0 0 3.266-1.313 5.316 
               5.316 0 0 0 1.62-3.255l1.127-10.331v-.158l.873-7.876a2.724 2.724 0 0 0-.038-.998z"/>
    </symbol>

    <!-- Іконка "Налаштування" - використовується для кнопки "Налаштування" -->
    <symbol id="icon-settings" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3"
            d="M16 20a4 4 0 1 0 0-8 4 4 0 0 0 0 8z"/>
    </symbol>

    <!-- Іконка "Видалити" (смітник) - використовується для кнопки "Видалити" -->
    <symbol id="icon-trash-04" viewBox="0 0 32 32">
      <path stroke-linecap="round" stroke-linejoin="round" stroke-width="3.6"
            d="M4 8h24m-2.667 0-.935 14.026c-.14 2.104-.21 3.156-.665 3.954a4.007 4.007 0 0 1-1.731 1.62"/>
    </symbol>

  </defs>
</svg> -->